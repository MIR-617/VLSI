interface operation;
  
  logic clk,reset;
  logic [3:0] out;
  
endinterface
