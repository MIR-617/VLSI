module andg(input_a,input_b,output_y);
input input_a,input_b;
output output_y;
assign output_y=input_a&input_b;
endmodule:andg
