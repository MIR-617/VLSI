// Code for xnor_gate  
module xnor_gate(
  input a,
  input b,
  output y
);
  xnor(y,a,b);
endmodule
