//code for and_gate
module and_gate(
  input a,
  input b,
  output y
);
  and(y,a,b);
endmodule
