module top_module( input in, output out );
    buf(out,in);

endmodule
