interface operation;
  
  logic clk,rst_n,d;
  logic q,qb;
  
endinterface
