// Code for xor_gate  level
module xor_gate(
  input a,
  input b,
  output y
);
  xor(y,a,b);
endmodule
