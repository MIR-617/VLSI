// Code for or_gate  
module or_gate(
  input a,
  input b,
  output y
);
  or(y,a,b);
endmodule
