module and_g(
  input a,
  input b,
  output y
);
  and(y,a,b);
endmodule
