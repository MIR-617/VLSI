class transaction;
  
  rand bit clk;
  bit reset;
  bit [3:0]out;
  
endclass
