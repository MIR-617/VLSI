// Code for not_gate  
module not_gate(
  input a,
  output y
);
  not(y,a);
endmodule
