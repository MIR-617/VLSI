class transaction;
  
   logic clk;
   logic rst_n;
   rand d;
   bit q;
   bit qb;
  
endclass
