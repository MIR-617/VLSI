interface and_if;
  logic a,b;
  logic y;
endinterface
